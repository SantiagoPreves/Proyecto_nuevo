-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition
-- Created on Mon Nov 06 16:16:05 2023

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY subgrupo_c IS
    PORT (
        clock : IN STD_LOGIC;
        reset : IN STD_LOGIC := '0';
        S : IN STD_LOGIC_VECTOR(1 DOWNTO 0) := "00";
        Mi : OUT STD_LOGIC;
        Md : OUT STD_LOGIC
    );
END subgrupo_c;

ARCHITECTURE BEHAVIOR OF subgrupo_c IS
    TYPE type_fstate IS (E0,E1,E2,E3);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,S)
    BEGIN
        IF (reset='0') THEN
            reg_fstate <= E0;
            Mi <= '0';
            Md <= '0';
        ELSE
            Mi <= '0';
            Md <= '0';
            CASE fstate IS
                WHEN E0 =>
                    IF ((S(1 DOWNTO 0) = "00")) THEN
                        reg_fstate <= E0;
                    ELSIF ((S(1 DOWNTO 0) = "11")) THEN
                        reg_fstate <= E1;
                    ELSIF ((S(1 DOWNTO 0) = "01")) THEN
                        reg_fstate <= E2;
                    ELSIF ((S(1 DOWNTO 0) = "10")) THEN
                        reg_fstate <= E3;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= E0;
                    END IF;

                    Md <= '1';

                    Mi <= '1';
                WHEN E1 =>
                    IF ((S(1 DOWNTO 0) = "00")) THEN
                        reg_fstate <= E0;
                    ELSIF ((S(1 DOWNTO 0) = "11")) THEN
                        reg_fstate <= E1;
                    ELSIF ((S(1 DOWNTO 0) = "01")) THEN
                        reg_fstate <= E2;
                    ELSIF ((S(1 DOWNTO 0) = "10")) THEN
                        reg_fstate <= E3;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= E1;
                    END IF;

                    Md <= '0';

                    Mi <= '0';
                WHEN E2 =>
                    IF ((S(1 DOWNTO 0) = "00")) THEN
                        reg_fstate <= E0;
                    ELSIF ((S(1 DOWNTO 0) = "11")) THEN
                        reg_fstate <= E1;
                    ELSIF ((S(1 DOWNTO 0) = "01")) THEN
                        reg_fstate <= E2;
                    ELSIF ((S(1 DOWNTO 0) = "10")) THEN
                        reg_fstate <= E3;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= E2;
                    END IF;

                    Md <= '1';

                    Mi <= '0';
                WHEN E3 =>
                    IF ((S(1 DOWNTO 0) = "00")) THEN
                        reg_fstate <= E0;
                    ELSIF ((S(1 DOWNTO 0) = "11")) THEN
                        reg_fstate <= E1;
                    ELSIF ((S(1 DOWNTO 0) = "01")) THEN
                        reg_fstate <= E2;
                    ELSIF ((S(1 DOWNTO 0) = "10")) THEN
                        reg_fstate <= E3;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= E3;
                    END IF;

                    Md <= '0';

                    Mi <= '1';
                WHEN OTHERS => 
                    Mi <= 'X';
                    Md <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
